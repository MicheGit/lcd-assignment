x1 >< x2: un? bool.end . x1 << true . 0 | x2 >> y: lin!bool.end . y << false . 0