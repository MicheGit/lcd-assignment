x >< y: lin? bool.end . x << true.0