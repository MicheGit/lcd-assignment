x1 >< x2: lin? bool.end . x1 << true . 0 | x3 >> y. 0